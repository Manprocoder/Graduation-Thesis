// system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module system (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] active_ascon_0_master_read_readdata;                         // mm_interconnect_0:active_ascon_0_Master_Read_readdata -> active_ascon_0:iReadData_Master_Read
	wire         active_ascon_0_master_read_waitrequest;                      // mm_interconnect_0:active_ascon_0_Master_Read_waitrequest -> active_ascon_0:iWait_Master_Read
	wire  [31:0] active_ascon_0_master_read_address;                          // active_ascon_0:oAddress_Master_Read -> mm_interconnect_0:active_ascon_0_Master_Read_address
	wire         active_ascon_0_master_read_read;                             // active_ascon_0:oRead_Master_Read -> mm_interconnect_0:active_ascon_0_Master_Read_read
	wire         active_ascon_0_master_read_readdatavalid;                    // mm_interconnect_0:active_ascon_0_Master_Read_readdatavalid -> active_ascon_0:iDataValid_Master_Read
	wire         active_ascon_0_master_write_waitrequest;                     // mm_interconnect_0:active_ascon_0_Master_Write_waitrequest -> active_ascon_0:iWait_Master_Write
	wire  [31:0] active_ascon_0_master_write_address;                         // active_ascon_0:oAddress_Master_Write -> mm_interconnect_0:active_ascon_0_Master_Write_address
	wire  [31:0] active_ascon_0_master_write_writedata;                       // active_ascon_0:oData_Master_Write -> mm_interconnect_0:active_ascon_0_Master_Write_writedata
	wire         active_ascon_0_master_write_write;                           // active_ascon_0:oWrite_Master_Write -> mm_interconnect_0:active_ascon_0_Master_Write_write
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [16:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [16:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_onchip_memory2_2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_2_s1_chipselect -> onchip_memory2_2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_2_s1_readdata;              // onchip_memory2_2:readdata -> mm_interconnect_0:onchip_memory2_2_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_2_s1_address;               // mm_interconnect_0:onchip_memory2_2_s1_address -> onchip_memory2_2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_2_s1_byteenable -> onchip_memory2_2:byteenable
	wire         mm_interconnect_0_onchip_memory2_2_s1_write;                 // mm_interconnect_0:onchip_memory2_2_s1_write -> onchip_memory2_2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_2_s1_writedata;             // mm_interconnect_0:onchip_memory2_2_s1_writedata -> onchip_memory2_2:writedata
	wire         mm_interconnect_0_onchip_memory2_2_s1_clken;                 // mm_interconnect_0:onchip_memory2_2_s1_clken -> onchip_memory2_2:clken
	wire         mm_interconnect_0_onchip_memory2_1_s1_chipselect;            // mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_readdata;              // onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_1_s1_address;               // mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_1_s1_byteenable;            // mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	wire         mm_interconnect_0_onchip_memory2_1_s1_write;                 // mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_writedata;             // mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	wire         mm_interconnect_0_onchip_memory2_1_s1_clken;                 // mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_active_ascon_0_control_slave_chipselect;   // mm_interconnect_0:active_ascon_0_control_slave_chipselect -> active_ascon_0:iChipSelect_Control
	wire  [31:0] mm_interconnect_0_active_ascon_0_control_slave_readdata;     // active_ascon_0:oData_Control -> mm_interconnect_0:active_ascon_0_control_slave_readdata
	wire   [1:0] mm_interconnect_0_active_ascon_0_control_slave_address;      // mm_interconnect_0:active_ascon_0_control_slave_address -> active_ascon_0:iAddress_Control
	wire         mm_interconnect_0_active_ascon_0_control_slave_read;         // mm_interconnect_0:active_ascon_0_control_slave_read -> active_ascon_0:iRead_Control
	wire         mm_interconnect_0_active_ascon_0_control_slave_write;        // mm_interconnect_0:active_ascon_0_control_slave_write -> active_ascon_0:iWrite_Control
	wire  [31:0] mm_interconnect_0_active_ascon_0_control_slave_writedata;    // mm_interconnect_0:active_ascon_0_control_slave_writedata -> active_ascon_0:iData_Control
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [active_ascon_0:iRstn, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:active_ascon_0_reset_sink_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, onchip_memory2_1:reset, onchip_memory2_2:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, onchip_memory2_1:reset_req, onchip_memory2_2:reset_req, rst_translator:reset_req_in]

	active_ascon #(
		.ROUNDS_PER_CYCLE0 (3),
		.ROUNDS_PER_CYCLE1 (2)
	) active_ascon_0 (
		.iClk                   (clk_clk),                                                   //    clock_sink.clk
		.iRstn                  (~rst_controller_reset_out_reset),                           //    reset_sink.reset_n
		.iChipSelect_Control    (mm_interconnect_0_active_ascon_0_control_slave_chipselect), // control_slave.chipselect
		.iWrite_Control         (mm_interconnect_0_active_ascon_0_control_slave_write),      //              .write
		.iRead_Control          (mm_interconnect_0_active_ascon_0_control_slave_read),       //              .read
		.iAddress_Control       (mm_interconnect_0_active_ascon_0_control_slave_address),    //              .address
		.iData_Control          (mm_interconnect_0_active_ascon_0_control_slave_writedata),  //              .writedata
		.oData_Control          (mm_interconnect_0_active_ascon_0_control_slave_readdata),   //              .readdata
		.oAddress_Master_Read   (active_ascon_0_master_read_address),                        //   Master_Read.address
		.oRead_Master_Read      (active_ascon_0_master_read_read),                           //              .read
		.iDataValid_Master_Read (active_ascon_0_master_read_readdatavalid),                  //              .readdatavalid
		.iReadData_Master_Read  (active_ascon_0_master_read_readdata),                       //              .readdata
		.iWait_Master_Read      (active_ascon_0_master_read_waitrequest),                    //              .waitrequest
		.oAddress_Master_Write  (active_ascon_0_master_write_address),                       //  Master_Write.address
		.oData_Master_Write     (active_ascon_0_master_write_writedata),                     //              .writedata
		.oWrite_Master_Write    (active_ascon_0_master_write_write),                         //              .write
		.iWait_Master_Write     (active_ascon_0_master_write_waitrequest)                    //              .waitrequest
	);

	system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	system_onchip_memory2_1 onchip_memory2_1 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	system_onchip_memory2_2 onchip_memory2_2 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                         (clk_clk),                                                     //                                       clock_clk.clk
		.active_ascon_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // active_ascon_0_reset_sink_reset_bridge_in_reset.reset
		.active_ascon_0_Master_Read_address                    (active_ascon_0_master_read_address),                          //                      active_ascon_0_Master_Read.address
		.active_ascon_0_Master_Read_waitrequest                (active_ascon_0_master_read_waitrequest),                      //                                                .waitrequest
		.active_ascon_0_Master_Read_read                       (active_ascon_0_master_read_read),                             //                                                .read
		.active_ascon_0_Master_Read_readdata                   (active_ascon_0_master_read_readdata),                         //                                                .readdata
		.active_ascon_0_Master_Read_readdatavalid              (active_ascon_0_master_read_readdatavalid),                    //                                                .readdatavalid
		.active_ascon_0_Master_Write_address                   (active_ascon_0_master_write_address),                         //                     active_ascon_0_Master_Write.address
		.active_ascon_0_Master_Write_waitrequest               (active_ascon_0_master_write_waitrequest),                     //                                                .waitrequest
		.active_ascon_0_Master_Write_write                     (active_ascon_0_master_write_write),                           //                                                .write
		.active_ascon_0_Master_Write_writedata                 (active_ascon_0_master_write_writedata),                       //                                                .writedata
		.nios2_gen2_0_data_master_address                      (nios2_gen2_0_data_master_address),                            //                        nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                  (nios2_gen2_0_data_master_waitrequest),                        //                                                .waitrequest
		.nios2_gen2_0_data_master_byteenable                   (nios2_gen2_0_data_master_byteenable),                         //                                                .byteenable
		.nios2_gen2_0_data_master_read                         (nios2_gen2_0_data_master_read),                               //                                                .read
		.nios2_gen2_0_data_master_readdata                     (nios2_gen2_0_data_master_readdata),                           //                                                .readdata
		.nios2_gen2_0_data_master_write                        (nios2_gen2_0_data_master_write),                              //                                                .write
		.nios2_gen2_0_data_master_writedata                    (nios2_gen2_0_data_master_writedata),                          //                                                .writedata
		.nios2_gen2_0_data_master_debugaccess                  (nios2_gen2_0_data_master_debugaccess),                        //                                                .debugaccess
		.nios2_gen2_0_instruction_master_address               (nios2_gen2_0_instruction_master_address),                     //                 nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest           (nios2_gen2_0_instruction_master_waitrequest),                 //                                                .waitrequest
		.nios2_gen2_0_instruction_master_read                  (nios2_gen2_0_instruction_master_read),                        //                                                .read
		.nios2_gen2_0_instruction_master_readdata              (nios2_gen2_0_instruction_master_readdata),                    //                                                .readdata
		.active_ascon_0_control_slave_address                  (mm_interconnect_0_active_ascon_0_control_slave_address),      //                    active_ascon_0_control_slave.address
		.active_ascon_0_control_slave_write                    (mm_interconnect_0_active_ascon_0_control_slave_write),        //                                                .write
		.active_ascon_0_control_slave_read                     (mm_interconnect_0_active_ascon_0_control_slave_read),         //                                                .read
		.active_ascon_0_control_slave_readdata                 (mm_interconnect_0_active_ascon_0_control_slave_readdata),     //                                                .readdata
		.active_ascon_0_control_slave_writedata                (mm_interconnect_0_active_ascon_0_control_slave_writedata),    //                                                .writedata
		.active_ascon_0_control_slave_chipselect               (mm_interconnect_0_active_ascon_0_control_slave_chipselect),   //                                                .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                   jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_0_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_0_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.nios2_gen2_0_debug_mem_slave_address                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //                    nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                                .write
		.nios2_gen2_0_debug_mem_slave_read                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                                .read
		.nios2_gen2_0_debug_mem_slave_readdata                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                                .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                                .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                                .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                                .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                                .debugaccess
		.onchip_memory2_0_s1_address                           (mm_interconnect_0_onchip_memory2_0_s1_address),               //                             onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                             (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                                .write
		.onchip_memory2_0_s1_readdata                          (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                                .readdata
		.onchip_memory2_0_s1_writedata                         (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                                .writedata
		.onchip_memory2_0_s1_byteenable                        (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                                .byteenable
		.onchip_memory2_0_s1_chipselect                        (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                                .chipselect
		.onchip_memory2_0_s1_clken                             (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                                .clken
		.onchip_memory2_1_s1_address                           (mm_interconnect_0_onchip_memory2_1_s1_address),               //                             onchip_memory2_1_s1.address
		.onchip_memory2_1_s1_write                             (mm_interconnect_0_onchip_memory2_1_s1_write),                 //                                                .write
		.onchip_memory2_1_s1_readdata                          (mm_interconnect_0_onchip_memory2_1_s1_readdata),              //                                                .readdata
		.onchip_memory2_1_s1_writedata                         (mm_interconnect_0_onchip_memory2_1_s1_writedata),             //                                                .writedata
		.onchip_memory2_1_s1_byteenable                        (mm_interconnect_0_onchip_memory2_1_s1_byteenable),            //                                                .byteenable
		.onchip_memory2_1_s1_chipselect                        (mm_interconnect_0_onchip_memory2_1_s1_chipselect),            //                                                .chipselect
		.onchip_memory2_1_s1_clken                             (mm_interconnect_0_onchip_memory2_1_s1_clken),                 //                                                .clken
		.onchip_memory2_2_s1_address                           (mm_interconnect_0_onchip_memory2_2_s1_address),               //                             onchip_memory2_2_s1.address
		.onchip_memory2_2_s1_write                             (mm_interconnect_0_onchip_memory2_2_s1_write),                 //                                                .write
		.onchip_memory2_2_s1_readdata                          (mm_interconnect_0_onchip_memory2_2_s1_readdata),              //                                                .readdata
		.onchip_memory2_2_s1_writedata                         (mm_interconnect_0_onchip_memory2_2_s1_writedata),             //                                                .writedata
		.onchip_memory2_2_s1_byteenable                        (mm_interconnect_0_onchip_memory2_2_s1_byteenable),            //                                                .byteenable
		.onchip_memory2_2_s1_chipselect                        (mm_interconnect_0_onchip_memory2_2_s1_chipselect),            //                                                .chipselect
		.onchip_memory2_2_s1_clken                             (mm_interconnect_0_onchip_memory2_2_s1_clken)                  //                                                .clken
	);

	system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
